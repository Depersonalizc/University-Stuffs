`timescale 1ns/1ps

module alu_test;

reg[31 : 0] i_datain, gr1, gr2;
wire[31 : 0] out, hi, lo;
wire zero, overflow, neg;

alu testalu(i_datain, gr1, gr2, out, hi, lo, zero, overflow, neg);

initial
begin
$display("instruction:op:fc:   gr1  :   gr2  :  srcA  :  srcB  :   out  :   hi   :   lo   :z:o:n:PCSrc:memW:regW:regD:mem2Reg:ALUctrl");
$monitor("   %h:%h:%h:%h:%h:%h:%h:%h:%h:%h:%h:%h:%h:  %h  :  %h :  %h :  %h:%h:%h",
        i_datain, testalu.opcode, testalu.funct, gr1, gr2, testalu.srcA, testalu.srcB, out, hi, lo, zero, overflow, neg, testalu.PCSrc, testalu.memWrite, testalu.memWrite, testalu.regDst,testalu.memToReg, testalu.ALUctrl);


#10 i_datain<=32'b00000010001100101000000000100001;	//	addu $s0, $s1, $s2
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00000010001100101000000000100010;	//	sub $s0, $s1, $s2
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00000010001100101000000000100011;	//	subu $s0, $s1, $s2
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00000010001100101000000000100100;	//	and $s0, $s1, $s2
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00000010001100101000000000100101;	//	or $s0, $s1, $s2
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00000010001100101000000000100111;	//	nor $s0, $s1, $s2
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00000001001010100100000000100110;	//  xor $t0, $t1, $t2
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00000001001010100000000000011010;	//	div $t1, $t2
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00000001100010100000000000011011;	//	divu $t4, $t2
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00000000000100011000001010000000;	//	sll $s0, $s1, 10
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00000000000100011000001010000010;	//	srl $s0, $s1, 10
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00000010011100011000000000000110;	//	srlv $s0, $s1, $s3
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00000000000100011000001010000011;	//	sra $s0, $s1, 10
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00000010011100011000000000000111;	//	srav $s0, $s1, $s3
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00000010001100111000000000101010;	//	slt $s0, $s1, $s3
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00000010001100111000000000101011;	//	sltu $s0, $s1, $s3
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00000001010010110000000000011000;	//	mult $t2, $t3
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00000001001010000000000000011001;	//	multu $t1, $t0
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00100110001100000000000001100100;	//	addiu $s0, $s1, 100
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00110010001100000000000001100100;	//	andi $s0, $s1, 100
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00110110001100000000000001100100;	//	ori $s0, $s1, 100
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00111010001100000000000001100100;	// 	xori $s0, $s1, 100
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00101010001100000000000001100100;	//	slti $s0, $s1, 100
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00101110001100000000000001100100;	//	sltiu $s0, $s1, 100
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00010010000100011111111111111000;	//	beq $s0, $s1, I
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00010110000100011111111111100100;	//	bne $s0, $s1, R
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b10001110001100000000000001100100;	//	lw $s0, 100($s1)
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b10101110001100000000000001100100;	//	sw $s0, 100($s1)
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00000001001010100100000000100000;	//	add $t0, $t1, $t2
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00100001001010001111111110000101;	//	addi $t0, $t1, -123
gr1<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00000001010010010100000000000100;	//	sllv $t0, $t1, $t2
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 i_datain<=32'b00000001001010100100000000100000;	//	add $t0, $t1, $t2 (overflow)
gr1<=32'b0101_1101_1101_1101_1101_1101_1101_1101;
gr2<=32'b0100_1101_1101_1101_1101_1101_1101_1101;

#10 $finish;
end
endmodule